CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 25 80 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
143654930 0
0
6 Title:
5 Name:
0
0
0
44
2 +V
167 1095 1087 0 1 3
0 16
0
0 0 53488 180
3 3S3
-11 -22 10 -14
3 ON1
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 1069 1086 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
9 CC 7-Seg~
183 1249 71 0 18 19
10 30 29 28 27 26 25 24 2 83
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP2
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3618 0 0
0
0
4 4511
219 1149 222 0 14 29
0 84 85 3 4 2 16 16 24 25
26 27 28 29 30
0
0 0 12528 0
4 4511
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
9 CC 7-Seg~
183 1313 71 0 18 19
10 37 36 35 34 33 32 31 2 86
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP1
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
9 CC 7-Seg~
183 1390 71 0 18 19
10 44 43 42 41 40 39 38 2 87
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP3
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7734 0 0
0
0
9 CC 7-Seg~
183 1455 71 0 18 19
10 51 50 49 48 47 46 45 2 88
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP4
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9914 0 0
0
0
9 CC 7-Seg~
183 1538 71 0 18 19
10 58 57 56 55 54 53 52 2 89
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP5
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3747 0 0
0
0
9 CC 7-Seg~
183 1598 71 0 18 19
10 65 64 63 62 61 60 59 2 90
1 1 1 1 1 1 0 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP6
27 -5 62 3
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3549 0 0
0
0
4 4511
219 1148 350 0 14 29
0 5 6 7 8 2 16 16 31 32
33 34 35 36 37
0
0 0 12528 0
4 4511
-14 -60 14 -52
3 U17
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
4 4511
219 1147 542 0 14 29
0 91 9 10 11 2 16 16 38 39
40 41 42 43 44
0
0 0 12528 0
4 4511
-14 -60 14 -52
3 U19
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
4 4511
219 1146 670 0 14 29
0 12 13 14 15 2 16 16 45 46
47 48 49 50 51
0
0 0 12528 0
4 4511
-14 -60 14 -52
3 U18
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
4 4511
219 1146 879 0 14 29
0 92 18 19 17 2 16 16 52 53
54 55 56 57 58
0
0 0 12528 0
4 4511
-14 -60 14 -52
3 U20
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
4 4511
219 1145 1007 0 20 29
0 20 21 22 23 2 16 16 59 60
61 62 63 64 65 0 0 0 0 0
1
0
0 0 12528 0
4 4511
-14 -60 14 -52
3 U21
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
7 Ground~
168 1682 129 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
10 2-In NAND~
219 525 1016 0 3 22
0 3 6 69
0
0 0 112 180
4 4011
-7 -24 21 -16
4 U16A
-11 -25 17 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 15 0
1 U
4718 0 0
0
0
9 2-In AND~
219 101 988 0 3 22
0 71 69 70
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U15A
18 -5 46 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 14 0
1 U
3874 0 0
0
0
10 4-In NAND~
219 174 1052 0 5 22
0 5 68 7 67 71
0
0 0 112 180
6 74LS20
-21 -28 21 -20
4 U14A
-11 -28 17 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 13 0
1 U
6671 0 0
0
0
6 JK RN~
219 615 895 0 6 22
0 66 4 66 69 93 3
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U13B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 12 0
1 U
3789 0 0
0
0
6 JK RN~
219 527 894 0 6 22
0 66 5 66 69 94 4
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U13A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 12 0
1 U
4871 0 0
0
0
6 JK RN~
219 438 894 0 6 22
0 66 6 66 70 95 5
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U12B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 11 0
1 U
3750 0 0
0
0
6 JK RN~
219 348 893 0 6 22
0 66 7 66 70 68 6
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U12A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 11 0
1 U
8778 0 0
0
0
6 JK RN~
219 259 892 0 6 22
0 66 8 66 70 96 7
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U11B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 10 0
1 U
538 0 0
0
0
6 JK RN~
219 168 892 0 6 22
0 66 9 66 70 67 8
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U11A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 10 0
1 U
6843 0 0
0
0
2 +V
167 83 173 0 1 3
0 66
0
0 0 53488 0
3 3S3
-11 -22 10 -14
2 ON
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3136 0 0
0
0
10 4-In NAND~
219 156 683 0 5 22
0 12 74 14 73 75
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U7B
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 6 0
1 U
5950 0 0
0
0
6 JK RN~
219 704 577 0 6 22
0 66 10 66 76 97 9
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U10B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 9 0
1 U
5670 0 0
0
0
6 JK RN~
219 611 577 0 6 22
0 66 11 66 76 98 10
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
4 U10A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 9 0
1 U
6828 0 0
0
0
6 JK RN~
219 522 577 0 6 22
0 66 12 66 76 72 11
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U9B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 8 0
1 U
6735 0 0
0
0
6 JK RN~
219 431 577 0 6 22
0 66 13 66 75 99 12
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U9A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 8 0
1 U
8365 0 0
0
0
6 JK RN~
219 341 577 0 6 22
0 66 14 66 75 74 13
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 7 0
1 U
4132 0 0
0
0
6 JK RN~
219 255 577 0 6 22
0 66 15 66 75 100 14
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U8A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 7 0
1 U
4551 0 0
0
0
6 JK RN~
219 165 576 0 6 22
0 66 18 66 75 73 15
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U5B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 4 0
1 U
3635 0 0
0
0
10 3-In NAND~
219 519 681 0 4 22
0 9 10 72 76
0
0 0 624 180
6 74LS10
-21 -28 21 -20
3 U6B
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 5 0
1 U
3973 0 0
0
0
10 4-In NAND~
219 154 365 0 5 22
0 20 79 22 78 80
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U7A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 -461928715
65 0 0 0 2 1 6 0
1 U
3851 0 0
0
0
10 3-In NAND~
219 517 363 0 4 22
0 18 19 77 81
0
0 0 624 180
6 74LS10
-21 -28 21 -20
3 U6A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
8383 0 0
0
0
6 JK RN~
219 163 258 0 6 22
0 66 82 66 80 78 23
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
9334 0 0
0
0
6 JK RN~
219 253 259 0 6 22
0 66 23 66 80 101 22
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
7471 0 0
0
0
6 JK RN~
219 339 259 0 6 22
0 66 22 66 80 79 21
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
3334 0 0
0
0
6 JK RN~
219 429 259 0 6 22
0 66 21 66 80 102 20
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3559 0 0
0
0
6 JK RN~
219 520 259 0 6 22
0 66 20 66 81 77 17
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 3 0
1 U
984 0 0
0
0
6 JK RN~
219 609 259 0 6 22
0 66 17 66 81 103 19
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U4B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 3 0
1 U
7557 0 0
0
0
6 JK RN~
219 702 259 0 6 22
0 66 19 66 81 104 18
0
0 0 4208 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 4 0
1 U
3146 0 0
0
0
7 Pulser~
4 31 243 0 10 12
0 105 106 82 107 0 0 2 2 1
7
0
0 0 4656 0
0
6 PULSER
-21 -28 21 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5687 0 0
0
0
188
0 3 3 0 0 12416 0 0 4 133 0 5
651 878
651 780
860 780
860 204
1117 204
0 4 4 0 0 12416 0 0 4 134 0 5
556 877
556 787
853 787
853 213
1117 213
0 1 5 0 0 12416 0 0 10 135 0 5
481 877
481 794
832 794
832 314
1116 314
0 2 6 0 0 12416 0 0 10 136 0 5
394 876
394 800
839 800
839 323
1116 323
0 3 7 0 0 8320 0 0 10 137 0 5
302 875
302 808
847 808
847 332
1116 332
0 4 8 0 0 8320 0 0 10 138 0 5
202 875
202 814
821 814
821 341
1116 341
2 0 9 0 0 8192 0 11 0 0 150 6
1115 515
1115 519
739 519
739 555
734 555
734 560
0 3 10 0 0 8320 0 0 11 162 0 5
642 560
642 526
1101 526
1101 524
1115 524
0 4 11 0 0 8320 0 0 11 163 0 3
557 560
557 533
1115 533
0 1 12 0 0 8320 0 0 12 164 0 5
460 560
460 541
820 541
820 634
1114 634
0 2 13 0 0 8320 0 0 12 165 0 5
377 560
377 533
841 533
841 643
1114 643
0 3 14 0 0 8320 0 0 12 166 0 5
286 560
286 541
826 541
826 652
1114 652
4 0 15 0 0 12416 0 12 0 0 167 5
1114 661
834 661
834 536
202 536
202 559
0 5 2 0 0 4096 0 0 12 31 0 2
1069 670
1108 670
0 5 2 0 0 4096 0 0 11 31 0 2
1069 542
1109 542
0 5 2 0 0 4096 0 0 10 31 0 2
1069 350
1110 350
0 7 16 0 0 4096 0 0 4 28 0 4
1095 241
1103 241
1103 240
1111 240
0 7 16 0 0 0 0 0 10 28 0 4
1095 369
1102 369
1102 368
1110 368
0 6 16 0 0 0 0 0 10 28 0 4
1095 360
1102 360
1102 359
1110 359
0 6 16 0 0 4096 0 0 11 28 0 2
1095 551
1109 551
0 7 16 0 0 0 0 0 11 28 0 2
1095 560
1109 560
0 6 16 0 0 0 0 0 12 28 0 4
1095 680
1100 680
1100 679
1108 679
0 7 16 0 0 0 0 0 12 28 0 2
1095 688
1108 688
0 7 16 0 0 0 0 0 13 28 0 2
1095 897
1108 897
0 6 16 0 0 0 0 0 13 28 0 2
1095 888
1108 888
0 7 16 0 0 0 0 0 14 28 0 2
1095 1025
1107 1025
0 6 16 0 0 0 0 0 14 28 0 4
1095 1017
1099 1017
1099 1016
1107 1016
1 6 16 0 0 4224 0 1 4 0 0 3
1095 1072
1095 231
1111 231
0 5 2 0 0 0 0 0 13 31 0 2
1069 879
1108 879
0 5 2 0 0 0 0 0 14 31 0 2
1069 1007
1107 1007
1 5 2 0 0 4224 0 2 4 0 0 3
1069 1080
1069 222
1111 222
4 0 17 0 0 8320 0 13 0 0 184 5
1114 870
813 870
813 222
560 222
560 242
0 2 18 0 0 12416 0 0 13 170 0 5
734 242
734 223
798 223
798 852
1114 852
0 3 19 0 0 12416 0 0 13 183 0 5
639 242
639 231
806 231
806 861
1114 861
0 1 20 0 0 12416 0 0 14 185 0 5
471 242
471 181
761 181
761 971
1113 971
0 2 21 0 0 12416 0 0 14 186 0 5
372 242
372 187
770 187
770 980
1113 980
0 3 22 0 0 12416 0 0 14 187 0 5
282 242
282 194
780 194
780 989
1113 989
0 4 23 0 0 12416 0 0 14 188 0 5
197 241
197 200
788 200
788 998
1113 998
8 7 24 0 0 8320 0 4 3 0 0 3
1181 240
1264 240
1264 107
9 6 25 0 0 8320 0 4 3 0 0 3
1181 231
1258 231
1258 107
10 5 26 0 0 8320 0 4 3 0 0 3
1181 222
1252 222
1252 107
11 4 27 0 0 8320 0 4 3 0 0 3
1181 213
1246 213
1246 107
12 3 28 0 0 8320 0 4 3 0 0 3
1181 204
1240 204
1240 107
13 2 29 0 0 8320 0 4 3 0 0 3
1181 195
1234 195
1234 107
14 1 30 0 0 8320 0 4 3 0 0 3
1181 186
1228 186
1228 107
8 7 31 0 0 8320 0 10 5 0 0 3
1180 368
1328 368
1328 107
9 6 32 0 0 8320 0 10 5 0 0 3
1180 359
1322 359
1322 107
10 5 33 0 0 8320 0 10 5 0 0 3
1180 350
1316 350
1316 107
11 4 34 0 0 8320 0 10 5 0 0 3
1180 341
1310 341
1310 107
12 3 35 0 0 8320 0 10 5 0 0 3
1180 332
1304 332
1304 107
13 2 36 0 0 8320 0 10 5 0 0 3
1180 323
1298 323
1298 107
14 1 37 0 0 8320 0 10 5 0 0 3
1180 314
1292 314
1292 107
0 8 2 0 0 0 0 0 5 86 0 2
1334 115
1334 107
8 7 38 0 0 8320 0 11 6 0 0 3
1179 560
1405 560
1405 107
9 6 39 0 0 8320 0 11 6 0 0 3
1179 551
1399 551
1399 107
10 5 40 0 0 8320 0 11 6 0 0 3
1179 542
1393 542
1393 107
11 4 41 0 0 8320 0 11 6 0 0 3
1179 533
1387 533
1387 107
12 3 42 0 0 8320 0 11 6 0 0 3
1179 524
1381 524
1381 107
13 2 43 0 0 8320 0 11 6 0 0 3
1179 515
1375 515
1375 107
14 1 44 0 0 8320 0 11 6 0 0 3
1179 506
1369 506
1369 107
0 8 2 0 0 0 0 0 6 86 0 3
1413 115
1413 107
1411 107
8 7 45 0 0 8320 0 12 7 0 0 3
1178 688
1470 688
1470 107
9 6 46 0 0 8320 0 12 7 0 0 3
1178 679
1464 679
1464 107
10 5 47 0 0 8320 0 12 7 0 0 3
1178 670
1458 670
1458 107
11 4 48 0 0 8320 0 12 7 0 0 3
1178 661
1452 661
1452 107
12 3 49 0 0 8320 0 12 7 0 0 3
1178 652
1446 652
1446 107
13 2 50 0 0 8320 0 12 7 0 0 3
1178 643
1440 643
1440 107
14 1 51 0 0 8320 0 12 7 0 0 3
1178 634
1434 634
1434 107
0 8 2 0 0 0 0 0 7 86 0 3
1478 115
1478 107
1476 107
8 7 52 0 0 8320 0 13 8 0 0 3
1178 897
1553 897
1553 107
9 6 53 0 0 8320 0 13 8 0 0 3
1178 888
1547 888
1547 107
10 5 54 0 0 8320 0 13 8 0 0 3
1178 879
1541 879
1541 107
11 4 55 0 0 8320 0 13 8 0 0 3
1178 870
1535 870
1535 107
12 3 56 0 0 8320 0 13 8 0 0 3
1178 861
1529 861
1529 107
13 2 57 0 0 8320 0 13 8 0 0 3
1178 852
1523 852
1523 107
14 1 58 0 0 8320 0 13 8 0 0 3
1178 843
1517 843
1517 107
0 8 2 0 0 0 0 0 8 86 0 3
1561 115
1561 107
1559 107
8 7 59 0 0 8320 0 14 9 0 0 3
1177 1025
1613 1025
1613 107
9 6 60 0 0 8320 0 14 9 0 0 3
1177 1016
1607 1016
1607 107
10 5 61 0 0 8320 0 14 9 0 0 3
1177 1007
1601 1007
1601 107
11 4 62 0 0 8320 0 14 9 0 0 3
1177 998
1595 998
1595 107
12 3 63 0 0 8320 0 14 9 0 0 3
1177 989
1589 989
1589 107
13 2 64 0 0 8320 0 14 9 0 0 3
1177 980
1583 980
1583 107
14 1 65 0 0 8320 0 14 9 0 0 3
1177 971
1577 971
1577 107
0 8 2 0 0 0 0 0 9 86 0 3
1624 115
1624 107
1619 107
1 8 2 0 0 0 0 15 3 0 0 4
1682 123
1682 115
1270 115
1270 107
0 1 66 0 0 8192 0 0 37 88 0 4
130 293
124 293
124 241
139 241
0 3 66 0 0 0 0 0 37 100 0 5
130 292
130 293
124 293
124 259
139 259
0 1 66 0 0 0 0 0 38 90 0 3
218 294
218 242
229 242
0 3 66 0 0 0 0 0 38 100 0 5
223 292
223 294
214 294
214 260
229 260
0 1 66 0 0 0 0 0 39 92 0 3
302 294
302 242
315 242
0 3 66 0 0 0 0 0 39 100 0 5
310 292
310 294
300 294
300 260
315 260
0 1 66 0 0 0 0 0 40 94 0 3
393 294
393 242
405 242
0 3 66 0 0 0 0 0 40 100 0 5
399 292
399 294
390 294
390 260
405 260
0 1 66 0 0 0 0 0 41 96 0 3
483 294
483 242
496 242
0 3 66 0 0 0 0 0 41 100 0 5
489 292
489 294
481 294
481 260
496 260
0 1 66 0 0 0 0 0 42 98 0 3
570 294
570 242
585 242
0 3 66 0 0 0 0 0 42 100 0 5
579 292
579 294
570 294
570 260
585 260
0 1 66 0 0 0 0 0 43 100 0 3
662 292
662 242
678 242
0 3 66 0 0 4096 0 0 43 126 0 4
83 292
663 292
663 260
678 260
0 1 66 0 0 0 0 0 33 102 0 3
126 612
126 559
141 559
0 3 66 0 0 0 0 0 33 114 0 3
126 612
126 577
141 577
0 1 66 0 0 0 0 0 32 104 0 3
216 612
216 560
231 560
0 3 66 0 0 0 0 0 32 114 0 4
222 612
216 612
216 578
231 578
0 1 66 0 0 0 0 0 31 106 0 3
302 612
302 560
317 560
0 3 66 0 0 0 0 0 31 114 0 4
312 612
302 612
302 578
317 578
0 1 66 0 0 0 0 0 30 108 0 3
393 612
393 560
407 560
0 3 66 0 0 0 0 0 30 114 0 4
402 612
392 612
392 578
407 578
0 1 66 0 0 0 0 0 29 110 0 3
483 612
483 560
498 560
0 3 66 0 0 0 0 0 29 114 0 3
483 612
483 578
498 578
0 1 66 0 0 0 0 0 28 112 0 3
574 612
574 560
587 560
0 3 66 0 0 0 0 0 28 114 0 4
584 612
572 612
572 578
587 578
0 1 66 0 0 0 0 0 27 114 0 3
665 612
665 560
680 560
0 3 66 0 0 4096 0 0 27 126 0 4
83 612
665 612
665 578
680 578
0 1 66 0 0 0 0 0 24 116 0 3
129 929
129 875
144 875
0 3 66 0 0 0 0 0 24 126 0 3
129 929
129 893
144 893
0 1 66 0 0 0 0 0 23 118 0 3
220 928
220 875
235 875
0 3 66 0 0 0 0 0 23 126 0 3
220 929
220 893
235 893
0 1 66 0 0 0 0 0 22 120 0 3
309 929
309 876
324 876
0 3 66 0 0 0 0 0 22 126 0 3
309 929
309 894
324 894
0 1 66 0 0 0 0 0 21 122 0 3
399 929
399 877
414 877
0 3 66 0 0 0 0 0 21 126 0 4
406 929
399 929
399 895
414 895
0 1 66 0 0 0 0 0 20 124 0 3
489 929
489 877
503 877
0 3 66 0 0 0 0 0 20 126 0 4
496 929
488 929
488 895
503 895
0 1 66 0 0 0 0 0 19 126 0 4
576 929
576 877
591 877
591 878
1 3 66 0 0 4224 0 25 19 0 0 5
83 182
83 929
576 929
576 896
591 896
0 2 9 0 0 8320 0 0 24 150 0 5
558 690
558 705
129 705
129 884
137 884
5 4 67 0 0 8320 0 24 18 0 0 4
198 893
208 893
208 1038
198 1038
0 3 7 0 0 0 0 0 18 137 0 3
295 875
295 1047
198 1047
5 2 68 0 0 12416 0 22 18 0 0 4
378 894
382 894
382 1056
198 1056
0 1 5 0 0 0 0 0 18 135 0 3
473 877
473 1065
198 1065
0 2 6 0 0 0 0 0 16 136 0 5
385 876
385 981
552 981
552 1007
549 1007
6 1 3 0 0 0 0 19 16 0 0 4
639 878
675 878
675 1025
549 1025
6 2 4 0 0 0 0 20 19 0 0 4
551 877
576 877
576 887
584 887
6 2 5 0 0 0 0 21 20 0 0 4
462 877
488 877
488 886
496 886
6 2 6 0 0 0 0 22 21 0 0 4
372 876
399 876
399 886
407 886
6 2 7 0 0 0 0 23 22 0 0 4
283 875
309 875
309 885
317 885
6 2 8 0 0 0 0 24 23 0 0 4
192 875
220 875
220 884
228 884
0 4 69 0 0 4096 0 0 20 140 0 2
527 934
527 925
0 4 69 0 0 8192 0 0 19 145 0 4
489 1016
489 934
615 934
615 926
0 4 70 0 0 4096 0 0 24 144 0 3
167 933
167 923
168 923
0 4 70 0 0 0 0 0 23 144 0 2
259 933
259 923
0 4 70 0 0 0 0 0 22 144 0 3
349 933
349 924
348 924
3 4 70 0 0 8320 0 17 21 0 0 4
100 964
100 933
438 933
438 925
3 2 69 0 0 4224 0 16 17 0 0 3
498 1016
109 1016
109 1009
5 1 71 0 0 4224 0 18 17 0 0 3
147 1052
91 1052
91 1009
0 2 18 0 0 0 0 0 33 170 0 5
556 372
556 388
126 388
126 568
134 568
5 3 72 0 0 8320 0 29 34 0 0 4
552 578
556 578
556 672
543 672
0 2 10 0 0 0 0 0 34 162 0 3
647 560
647 681
543 681
6 1 9 0 0 0 0 27 34 0 0 4
728 560
738 560
738 690
543 690
5 4 73 0 0 8320 0 33 26 0 0 4
195 577
199 577
199 669
180 669
0 3 14 0 0 0 0 0 26 166 0 3
290 560
290 678
180 678
5 2 74 0 0 12416 0 31 26 0 0 4
371 578
375 578
375 687
180 687
0 1 12 0 0 0 0 0 26 164 0 3
464 560
464 696
180 696
0 4 75 0 0 4096 0 0 31 161 0 3
342 616
342 608
341 608
0 4 75 0 0 0 0 0 32 161 0 3
256 616
256 608
255 608
0 4 75 0 0 4096 0 0 33 161 0 3
166 616
166 607
165 607
0 4 76 0 0 4096 0 0 29 160 0 2
522 616
522 608
4 0 76 0 0 0 0 28 0 0 160 2
611 608
611 616
4 4 76 0 0 12416 0 34 27 0 0 5
492 681
490 681
490 616
704 616
704 608
5 4 75 0 0 12416 0 26 30 0 0 5
129 683
127 683
127 616
431 616
431 608
6 2 10 0 0 0 0 28 27 0 0 4
635 560
665 560
665 569
673 569
6 2 11 0 0 0 0 29 28 0 0 4
546 560
572 560
572 569
580 569
6 2 12 0 0 0 0 30 29 0 0 4
455 560
483 560
483 569
491 569
6 2 13 0 0 0 0 31 30 0 0 4
365 560
392 560
392 569
400 569
6 2 14 0 0 0 0 32 31 0 0 4
279 560
302 560
302 569
310 569
6 2 15 0 0 0 0 33 32 0 0 4
189 559
216 559
216 569
224 569
5 3 77 0 0 8320 0 41 36 0 0 4
550 260
554 260
554 354
541 354
0 2 19 0 0 0 0 0 36 183 0 3
645 242
645 363
541 363
6 1 18 0 0 0 0 43 36 0 0 4
726 242
736 242
736 372
541 372
5 4 78 0 0 8320 0 37 35 0 0 4
193 259
197 259
197 351
178 351
0 3 22 0 0 0 0 0 35 187 0 3
288 242
288 360
178 360
5 2 79 0 0 12416 0 39 35 0 0 4
369 260
373 260
373 369
178 369
0 1 20 0 0 0 0 0 35 185 0 3
462 242
462 378
178 378
0 4 80 0 0 4096 0 0 39 181 0 3
340 298
340 290
339 290
0 4 80 0 0 0 0 0 38 181 0 3
254 298
254 290
253 290
0 4 80 0 0 4096 0 0 37 181 0 3
164 298
164 289
163 289
0 4 81 0 0 4096 0 0 41 180 0 2
520 298
520 290
4 0 81 0 0 0 0 42 0 0 180 2
609 290
609 298
4 4 81 0 0 12416 0 36 43 0 0 5
490 363
488 363
488 298
702 298
702 290
5 4 80 0 0 12416 0 35 40 0 0 5
127 365
125 365
125 298
429 298
429 290
3 2 82 0 0 4224 0 44 37 0 0 4
55 234
124 234
124 250
132 250
6 2 19 0 0 0 0 42 43 0 0 4
633 242
663 242
663 251
671 251
6 2 17 0 0 0 0 41 42 0 0 4
544 242
570 242
570 251
578 251
6 2 20 0 0 0 0 40 41 0 0 4
453 242
481 242
481 251
489 251
6 2 21 0 0 0 0 39 40 0 0 4
363 242
390 242
390 251
398 251
6 2 22 0 0 0 0 38 39 0 0 4
277 242
300 242
300 251
308 251
6 2 23 0 0 0 0 37 38 0 0 4
187 241
214 241
214 251
222 251
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
85 150 241 173
98 160 246 175
21 Mantem J e K sempre 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
1064 137 1205 160
1077 147 1210 162
19 DECODIFICADOR HORAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
1103 452 1259 475
1116 462 1264 477
21 DECODIFICADOR MINUTOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1100 789 1262 812
1112 799 1266 814
22 DECODIFICADOR SEGUNDOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
349 482 406 505
361 492 410 507
7 MINUTOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
354 760 402 784
364 768 404 784
5 HORAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1387 6 1444 29
1399 16 1448 31
7 MINUTOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1257 9 1305 33
1267 17 1307 33
5 HORAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
367 135 431 158
380 145 436 160
8 SEGUNDOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1527 4 1591 27
1540 14 1596 29
8 SEGUNDOS
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
